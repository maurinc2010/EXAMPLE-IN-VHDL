library verilog;
use verilog.vl_types.all;
entity SEMAFORO_vlg_vec_tst is
end SEMAFORO_vlg_vec_tst;
