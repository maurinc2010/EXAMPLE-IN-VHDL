library verilog;
use verilog.vl_types.all;
entity TECLADO_vlg_vec_tst is
end TECLADO_vlg_vec_tst;
